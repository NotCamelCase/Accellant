`ifndef __CONFIG_SVH__
`define __CONFIG_SVH__

// Toggle forwarding result from WB stage to save one cycle during Dispatch
parameter   ENABLE_BYPASS_WB    = 1'b0;

`endif